library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity BN_to_BCD is
    Port (
        BN 		: in  STD_LOGIC_VECTOR(5 downto 0);  
        Dig_1  : out STD_LOGIC_VECTOR(3 downto 0); 
        Dig_2  : out STD_LOGIC_VECTOR(3 downto 0)  
    );
end BN_to_BCD;

architecture Behavioral of BN_to_BCD is
begin
    process(BN)
    begin

        case BN is
            when "000000" =>
                -- Decimal 0
                Dig_1 <= "0000";
                Dig_2 <= "0000";
            when "000001" =>
                -- Decimal 1
                Dig_1 <= "0000";
                Dig_2 <= "0001";
            when "000010" =>
                -- Decimal 2
                Dig_1 <= "0000";
                Dig_2 <= "0010";
            when "000011" =>
                -- Decimal 3
                Dig_1 <= "0000";
                Dig_2 <= "0011";
            when "000100" =>
                -- Decimal 4
                Dig_1 <= "0000";
                Dig_2 <= "0100";
            when "000101" =>
                -- Decimal 5
                Dig_1 <= "0000";
                Dig_2 <= "0101";
            when "000110" =>
                -- Decimal 6
                Dig_1 <= "0000";
                Dig_2 <= "0110";
            when "000111" =>
                -- Decimal 7
                Dig_1 <= "0000";
                Dig_2 <= "0111";
            when "001000" =>
                -- Decimal 8
                Dig_1 <= "0000";
                Dig_2 <= "1000";
            when "001001" =>
                -- Decimal 9
                Dig_1 <= "0000";
                Dig_2 <= "1001";
            when "001010" => -- Decimal 10
                Dig_1 <= "0001";
                Dig_2 <= "0000";
            when "001011" =>
                -- Decimal 11
                Dig_1 <= "0001";
                Dig_2 <= "0001";
            when "001100" =>
                -- Decimal 12
                Dig_1 <= "0001";
                Dig_2 <= "0010";
            when "001101" =>
                -- Decimal 13
                Dig_1 <= "0001";
                Dig_2 <= "0011";
            when "001110" =>
                -- Decimal 14
                Dig_1 <= "0001";
                Dig_2 <= "0100";
            when "001111" =>
                -- Decimal 15
                Dig_1 <= "0001";
                Dig_2 <= "0101";
            when "010000" =>
                -- Decimal 16
                Dig_1 <= "0001";
                Dig_2 <= "0110";
            when "010001" =>
                -- Decimal 17
                Dig_1 <= "0001";
                Dig_2 <= "0111";
            when "010010" =>
                -- Decimal 18
                Dig_1 <= "0001";
                Dig_2 <= "1000";
            when "010011" =>
                -- Decimal 19
                Dig_1 <= "0001";
                Dig_2 <= "1001";
            when "010100" => -- Decimal 20
                Dig_1 <= "0010";
                Dig_2 <= "0000";
            when "010101" =>
                -- Decimal 21
                Dig_1 <= "0010";
                Dig_2 <= "0001";
            when "010110" =>
                -- Decimal 22
                Dig_1 <= "0010";
                Dig_2 <= "0010";
            when "010111" =>
                -- Decimal 23
                Dig_1 <= "0010";
                Dig_2 <= "0011";
            when "011000" =>
                -- Decimal 24
                Dig_1 <= "0010";
                Dig_2 <= "0100";
            when "011001" =>
                -- Decimal 25
                Dig_1 <= "0010";
                Dig_2 <= "0101";
            when "011010" =>
                -- Decimal 26
                Dig_1 <= "0010";
                Dig_2 <= "0110";
            when "011011" =>
                -- Decimal 27
                Dig_1 <= "0010";
                Dig_2 <= "0111";
            when "011100" =>
                -- Decimal 28
                Dig_1 <= "0010";
                Dig_2 <= "1000";
            when "011101" =>
                -- Decimal 29
                Dig_1 <= "0010";
                Dig_2 <= "1001";
            when "011110" =>
                -- Decimal 30
                Dig_1 <= "0011";
                Dig_2 <= "0000";
            when "011111" =>
                -- Decimal 31
                Dig_1 <= "0011";
                Dig_2 <= "0001";
            when "100000" =>
                -- Decimal 32
                Dig_1 <= "0011";
                Dig_2 <= "0010";
            when "100001" =>
                -- Decimal 33
                Dig_1 <= "0011";
                Dig_2 <= "0011";
            when "100010" =>
                -- Decimal 34
                Dig_1 <= "0011";
                Dig_2 <= "0100";
            when "100011" =>
                -- Decimal 35
                Dig_1 <= "0011";
                Dig_2 <= "0101";
            when "100100" =>
                -- Decimal 36
                Dig_1 <= "0011";
                Dig_2 <= "0110";
            when "100101" =>
                -- Decimal 37
                Dig_1 <= "0011";
                Dig_2 <= "0111";
            when "100110" =>
                -- Decimal 38
                Dig_1 <= "0011";
                Dig_2 <= "1000";
            when "100111" =>
                -- Decimal 39
                Dig_1 <= "0011";
                Dig_2 <= "1001";
            when "101000" =>
                -- Decimal 40
                Dig_1 <= "0100";
                Dig_2 <= "0000";
            when "101001" =>
                -- Decimal 41
                Dig_1 <= "0100";
                Dig_2 <= "0001";
            when "101010" =>
                -- Decimal 42
                Dig_1 <= "0100";
                Dig_2 <= "0010";
            when "101011" =>
                -- Decimal 43
                Dig_1 <= "0100";
                Dig_2 <= "0011";
            when "101100" =>
                -- Decimal 44
                Dig_1 <= "0100";
                Dig_2 <= "0100";
            when "101101" =>
                -- Decimal 45
                Dig_1 <= "0100";
                Dig_2 <= "0101";
            when "101110" =>
                -- Decimal 46
                Dig_1 <= "0100";
                Dig_2 <= "0110";
            when "101111" =>
                -- Decimal 47
                Dig_1 <= "0100";
                Dig_2 <= "0111";
            when "110000" =>
                -- Decimal 48
                Dig_1 <= "0100";
                Dig_2 <= "1000";
            when "110001" =>
                -- Decimal 49
                Dig_1 <= "0100";
                Dig_2 <= "1001";
            when "110010" =>
                -- Decimal 50
                Dig_1 <= "0101";
                Dig_2 <= "0000";
            when "110011" =>
                -- Decimal 51
                Dig_1 <= "0101";
                Dig_2 <= "0001";
            when "110100" =>
                -- Decimal 52
                Dig_1 <= "0101";
                Dig_2 <= "0010";
            when "110101" =>
                -- Decimal 53
                Dig_1 <= "0101";
                Dig_2 <= "0011";
            when "110110" =>
                -- Decimal 54
                Dig_1 <= "0101";
                Dig_2 <= "0100";
            when "110111" =>
                -- Decimal 55
                Dig_1 <= "0101";
                Dig_2 <= "0101";
            when "111000" =>
                -- Decimal 56
                Dig_1 <= "0101";
                Dig_2 <= "0110";
            when "111001" =>
                -- Decimal 57
                Dig_1 <= "0101";
                Dig_2 <= "0111";
            when "111010" =>
                -- Decimal 58
                Dig_1 <= "0101";
                Dig_2 <= "1000";
            when "111011" =>
                -- Decimal 59
                Dig_1 <= "0101";
                Dig_2 <= "1001";
            when "111100" =>
                -- Decimal 60
                Dig_1 <= "0110";
                Dig_2 <= "0000";
            when "111101" =>
                -- Decimal 61
                Dig_1 <= "0110";
                Dig_2 <= "0001";
            when "111110" =>
                -- Decimal 62
                Dig_1 <= "0110";
                Dig_2 <= "0010";
            when "111111" =>
                -- Decimal 63
                Dig_1 <= "0110";
                Dig_2 <= "0011";

            when others =>
                Dig_1 <= (others => '0');
                Dig_2 <= (others => '0');
        end case;
    end process;
end Behavioral;
